// signle-bit signal state detection
$rose(); $fell(); $stable();


// Input generation
array_1.randomize(); 
